//-----------------------------------------------------------------------------
// system_axi_perf_mon_0_wrapper.v
//-----------------------------------------------------------------------------

(* x_core_info = "axi_perf_mon_v3_00_a" *)
module system_axi_perf_mon_0_wrapper
  (
    S_AXI_ACLK,
    S_AXI_ARESETN,
    S_AXI_AWADDR,
    S_AXI_AWVALID,
    S_AXI_AWREADY,
    S_AXI_WDATA,
    S_AXI_WSTRB,
    S_AXI_WVALID,
    S_AXI_WREADY,
    S_AXI_BRESP,
    S_AXI_BVALID,
    S_AXI_BREADY,
    S_AXI_ARADDR,
    S_AXI_ARVALID,
    S_AXI_ARREADY,
    S_AXI_RDATA,
    S_AXI_RRESP,
    S_AXI_RVALID,
    S_AXI_RREADY,
    SLOT_0_AXI_ACLK,
    SLOT_0_AXI_ARESETN,
    SLOT_0_AXI_AWID,
    SLOT_0_AXI_AWADDR,
    SLOT_0_AXI_AWLEN,
    SLOT_0_AXI_AWPROT,
    SLOT_0_AXI_AWSIZE,
    SLOT_0_AXI_AWBURST,
    SLOT_0_AXI_AWCACHE,
    SLOT_0_AXI_AWLOCK,
    SLOT_0_AXI_AWVALID,
    SLOT_0_AXI_AWREADY,
    SLOT_0_AXI_WDATA,
    SLOT_0_AXI_WSTRB,
    SLOT_0_AXI_WLAST,
    SLOT_0_AXI_WVALID,
    SLOT_0_AXI_WREADY,
    SLOT_0_AXI_BID,
    SLOT_0_AXI_BRESP,
    SLOT_0_AXI_BVALID,
    SLOT_0_AXI_BREADY,
    SLOT_0_AXI_ARID,
    SLOT_0_AXI_ARADDR,
    SLOT_0_AXI_ARLEN,
    SLOT_0_AXI_ARSIZE,
    SLOT_0_AXI_ARBURST,
    SLOT_0_AXI_ARPROT,
    SLOT_0_AXI_ARCACHE,
    SLOT_0_AXI_ARLOCK,
    SLOT_0_AXI_ARVALID,
    SLOT_0_AXI_ARREADY,
    SLOT_0_AXI_RID,
    SLOT_0_AXI_RDATA,
    SLOT_0_AXI_RRESP,
    SLOT_0_AXI_RLAST,
    SLOT_0_AXI_RVALID,
    SLOT_0_AXI_RREADY,
    SLOT_0_AXIS_ACLK,
    SLOT_0_AXIS_ARESETN,
    SLOT_0_AXIS_TVALID,
    SLOT_0_AXIS_TREADY,
    SLOT_0_AXIS_TDATA,
    SLOT_0_AXIS_TSTRB,
    SLOT_0_AXIS_TKEEP,
    SLOT_0_AXIS_TLAST,
    SLOT_0_AXIS_TID,
    SLOT_0_AXIS_TDEST,
    SLOT_0_AXIS_TUSER,
    SLOT_1_AXI_ACLK,
    SLOT_1_AXI_ARESETN,
    SLOT_1_AXI_AWID,
    SLOT_1_AXI_AWADDR,
    SLOT_1_AXI_AWLEN,
    SLOT_1_AXI_AWPROT,
    SLOT_1_AXI_AWSIZE,
    SLOT_1_AXI_AWBURST,
    SLOT_1_AXI_AWCACHE,
    SLOT_1_AXI_AWLOCK,
    SLOT_1_AXI_AWVALID,
    SLOT_1_AXI_AWREADY,
    SLOT_1_AXI_WDATA,
    SLOT_1_AXI_WSTRB,
    SLOT_1_AXI_WLAST,
    SLOT_1_AXI_WVALID,
    SLOT_1_AXI_WREADY,
    SLOT_1_AXI_BID,
    SLOT_1_AXI_BRESP,
    SLOT_1_AXI_BVALID,
    SLOT_1_AXI_BREADY,
    SLOT_1_AXI_ARID,
    SLOT_1_AXI_ARADDR,
    SLOT_1_AXI_ARLEN,
    SLOT_1_AXI_ARSIZE,
    SLOT_1_AXI_ARBURST,
    SLOT_1_AXI_ARPROT,
    SLOT_1_AXI_ARCACHE,
    SLOT_1_AXI_ARLOCK,
    SLOT_1_AXI_ARVALID,
    SLOT_1_AXI_ARREADY,
    SLOT_1_AXI_RID,
    SLOT_1_AXI_RDATA,
    SLOT_1_AXI_RRESP,
    SLOT_1_AXI_RLAST,
    SLOT_1_AXI_RVALID,
    SLOT_1_AXI_RREADY,
    SLOT_1_AXIS_ACLK,
    SLOT_1_AXIS_ARESETN,
    SLOT_1_AXIS_TVALID,
    SLOT_1_AXIS_TREADY,
    SLOT_1_AXIS_TDATA,
    SLOT_1_AXIS_TSTRB,
    SLOT_1_AXIS_TKEEP,
    SLOT_1_AXIS_TLAST,
    SLOT_1_AXIS_TID,
    SLOT_1_AXIS_TDEST,
    SLOT_1_AXIS_TUSER,
    SLOT_2_AXI_ACLK,
    SLOT_2_AXI_ARESETN,
    SLOT_2_AXI_AWID,
    SLOT_2_AXI_AWADDR,
    SLOT_2_AXI_AWLEN,
    SLOT_2_AXI_AWPROT,
    SLOT_2_AXI_AWSIZE,
    SLOT_2_AXI_AWBURST,
    SLOT_2_AXI_AWCACHE,
    SLOT_2_AXI_AWLOCK,
    SLOT_2_AXI_AWVALID,
    SLOT_2_AXI_AWREADY,
    SLOT_2_AXI_WDATA,
    SLOT_2_AXI_WSTRB,
    SLOT_2_AXI_WLAST,
    SLOT_2_AXI_WVALID,
    SLOT_2_AXI_WREADY,
    SLOT_2_AXI_BID,
    SLOT_2_AXI_BRESP,
    SLOT_2_AXI_BVALID,
    SLOT_2_AXI_BREADY,
    SLOT_2_AXI_ARID,
    SLOT_2_AXI_ARADDR,
    SLOT_2_AXI_ARLEN,
    SLOT_2_AXI_ARSIZE,
    SLOT_2_AXI_ARBURST,
    SLOT_2_AXI_ARPROT,
    SLOT_2_AXI_ARCACHE,
    SLOT_2_AXI_ARLOCK,
    SLOT_2_AXI_ARVALID,
    SLOT_2_AXI_ARREADY,
    SLOT_2_AXI_RID,
    SLOT_2_AXI_RDATA,
    SLOT_2_AXI_RRESP,
    SLOT_2_AXI_RLAST,
    SLOT_2_AXI_RVALID,
    SLOT_2_AXI_RREADY,
    SLOT_2_AXIS_ACLK,
    SLOT_2_AXIS_ARESETN,
    SLOT_2_AXIS_TVALID,
    SLOT_2_AXIS_TREADY,
    SLOT_2_AXIS_TDATA,
    SLOT_2_AXIS_TSTRB,
    SLOT_2_AXIS_TKEEP,
    SLOT_2_AXIS_TLAST,
    SLOT_2_AXIS_TID,
    SLOT_2_AXIS_TDEST,
    SLOT_2_AXIS_TUSER,
    SLOT_3_AXI_ACLK,
    SLOT_3_AXI_ARESETN,
    SLOT_3_AXI_AWID,
    SLOT_3_AXI_AWADDR,
    SLOT_3_AXI_AWLEN,
    SLOT_3_AXI_AWPROT,
    SLOT_3_AXI_AWSIZE,
    SLOT_3_AXI_AWBURST,
    SLOT_3_AXI_AWCACHE,
    SLOT_3_AXI_AWLOCK,
    SLOT_3_AXI_AWVALID,
    SLOT_3_AXI_AWREADY,
    SLOT_3_AXI_WDATA,
    SLOT_3_AXI_WSTRB,
    SLOT_3_AXI_WLAST,
    SLOT_3_AXI_WVALID,
    SLOT_3_AXI_WREADY,
    SLOT_3_AXI_BID,
    SLOT_3_AXI_BRESP,
    SLOT_3_AXI_BVALID,
    SLOT_3_AXI_BREADY,
    SLOT_3_AXI_ARID,
    SLOT_3_AXI_ARADDR,
    SLOT_3_AXI_ARLEN,
    SLOT_3_AXI_ARSIZE,
    SLOT_3_AXI_ARBURST,
    SLOT_3_AXI_ARPROT,
    SLOT_3_AXI_ARCACHE,
    SLOT_3_AXI_ARLOCK,
    SLOT_3_AXI_ARVALID,
    SLOT_3_AXI_ARREADY,
    SLOT_3_AXI_RID,
    SLOT_3_AXI_RDATA,
    SLOT_3_AXI_RRESP,
    SLOT_3_AXI_RLAST,
    SLOT_3_AXI_RVALID,
    SLOT_3_AXI_RREADY,
    SLOT_3_AXIS_ACLK,
    SLOT_3_AXIS_ARESETN,
    SLOT_3_AXIS_TVALID,
    SLOT_3_AXIS_TREADY,
    SLOT_3_AXIS_TDATA,
    SLOT_3_AXIS_TSTRB,
    SLOT_3_AXIS_TKEEP,
    SLOT_3_AXIS_TLAST,
    SLOT_3_AXIS_TID,
    SLOT_3_AXIS_TDEST,
    SLOT_3_AXIS_TUSER,
    SLOT_4_AXI_ACLK,
    SLOT_4_AXI_ARESETN,
    SLOT_4_AXI_AWID,
    SLOT_4_AXI_AWADDR,
    SLOT_4_AXI_AWLEN,
    SLOT_4_AXI_AWPROT,
    SLOT_4_AXI_AWSIZE,
    SLOT_4_AXI_AWBURST,
    SLOT_4_AXI_AWCACHE,
    SLOT_4_AXI_AWLOCK,
    SLOT_4_AXI_AWVALID,
    SLOT_4_AXI_AWREADY,
    SLOT_4_AXI_WDATA,
    SLOT_4_AXI_WSTRB,
    SLOT_4_AXI_WLAST,
    SLOT_4_AXI_WVALID,
    SLOT_4_AXI_WREADY,
    SLOT_4_AXI_BID,
    SLOT_4_AXI_BRESP,
    SLOT_4_AXI_BVALID,
    SLOT_4_AXI_BREADY,
    SLOT_4_AXI_ARID,
    SLOT_4_AXI_ARADDR,
    SLOT_4_AXI_ARLEN,
    SLOT_4_AXI_ARSIZE,
    SLOT_4_AXI_ARBURST,
    SLOT_4_AXI_ARPROT,
    SLOT_4_AXI_ARCACHE,
    SLOT_4_AXI_ARLOCK,
    SLOT_4_AXI_ARVALID,
    SLOT_4_AXI_ARREADY,
    SLOT_4_AXI_RID,
    SLOT_4_AXI_RDATA,
    SLOT_4_AXI_RRESP,
    SLOT_4_AXI_RLAST,
    SLOT_4_AXI_RVALID,
    SLOT_4_AXI_RREADY,
    SLOT_4_AXIS_ACLK,
    SLOT_4_AXIS_ARESETN,
    SLOT_4_AXIS_TVALID,
    SLOT_4_AXIS_TREADY,
    SLOT_4_AXIS_TDATA,
    SLOT_4_AXIS_TSTRB,
    SLOT_4_AXIS_TKEEP,
    SLOT_4_AXIS_TLAST,
    SLOT_4_AXIS_TID,
    SLOT_4_AXIS_TDEST,
    SLOT_4_AXIS_TUSER,
    SLOT_5_AXI_ACLK,
    SLOT_5_AXI_ARESETN,
    SLOT_5_AXI_AWID,
    SLOT_5_AXI_AWADDR,
    SLOT_5_AXI_AWLEN,
    SLOT_5_AXI_AWPROT,
    SLOT_5_AXI_AWSIZE,
    SLOT_5_AXI_AWBURST,
    SLOT_5_AXI_AWCACHE,
    SLOT_5_AXI_AWLOCK,
    SLOT_5_AXI_AWVALID,
    SLOT_5_AXI_AWREADY,
    SLOT_5_AXI_WDATA,
    SLOT_5_AXI_WSTRB,
    SLOT_5_AXI_WLAST,
    SLOT_5_AXI_WVALID,
    SLOT_5_AXI_WREADY,
    SLOT_5_AXI_BID,
    SLOT_5_AXI_BRESP,
    SLOT_5_AXI_BVALID,
    SLOT_5_AXI_BREADY,
    SLOT_5_AXI_ARID,
    SLOT_5_AXI_ARADDR,
    SLOT_5_AXI_ARLEN,
    SLOT_5_AXI_ARSIZE,
    SLOT_5_AXI_ARBURST,
    SLOT_5_AXI_ARPROT,
    SLOT_5_AXI_ARCACHE,
    SLOT_5_AXI_ARLOCK,
    SLOT_5_AXI_ARVALID,
    SLOT_5_AXI_ARREADY,
    SLOT_5_AXI_RID,
    SLOT_5_AXI_RDATA,
    SLOT_5_AXI_RRESP,
    SLOT_5_AXI_RLAST,
    SLOT_5_AXI_RVALID,
    SLOT_5_AXI_RREADY,
    SLOT_5_AXIS_ACLK,
    SLOT_5_AXIS_ARESETN,
    SLOT_5_AXIS_TVALID,
    SLOT_5_AXIS_TREADY,
    SLOT_5_AXIS_TDATA,
    SLOT_5_AXIS_TSTRB,
    SLOT_5_AXIS_TKEEP,
    SLOT_5_AXIS_TLAST,
    SLOT_5_AXIS_TID,
    SLOT_5_AXIS_TDEST,
    SLOT_5_AXIS_TUSER,
    SLOT_6_AXI_ACLK,
    SLOT_6_AXI_ARESETN,
    SLOT_6_AXI_AWID,
    SLOT_6_AXI_AWADDR,
    SLOT_6_AXI_AWLEN,
    SLOT_6_AXI_AWPROT,
    SLOT_6_AXI_AWSIZE,
    SLOT_6_AXI_AWBURST,
    SLOT_6_AXI_AWCACHE,
    SLOT_6_AXI_AWLOCK,
    SLOT_6_AXI_AWVALID,
    SLOT_6_AXI_AWREADY,
    SLOT_6_AXI_WDATA,
    SLOT_6_AXI_WSTRB,
    SLOT_6_AXI_WLAST,
    SLOT_6_AXI_WVALID,
    SLOT_6_AXI_WREADY,
    SLOT_6_AXI_BID,
    SLOT_6_AXI_BRESP,
    SLOT_6_AXI_BVALID,
    SLOT_6_AXI_BREADY,
    SLOT_6_AXI_ARID,
    SLOT_6_AXI_ARADDR,
    SLOT_6_AXI_ARLEN,
    SLOT_6_AXI_ARSIZE,
    SLOT_6_AXI_ARBURST,
    SLOT_6_AXI_ARPROT,
    SLOT_6_AXI_ARCACHE,
    SLOT_6_AXI_ARLOCK,
    SLOT_6_AXI_ARVALID,
    SLOT_6_AXI_ARREADY,
    SLOT_6_AXI_RID,
    SLOT_6_AXI_RDATA,
    SLOT_6_AXI_RRESP,
    SLOT_6_AXI_RLAST,
    SLOT_6_AXI_RVALID,
    SLOT_6_AXI_RREADY,
    SLOT_6_AXIS_ACLK,
    SLOT_6_AXIS_ARESETN,
    SLOT_6_AXIS_TVALID,
    SLOT_6_AXIS_TREADY,
    SLOT_6_AXIS_TDATA,
    SLOT_6_AXIS_TSTRB,
    SLOT_6_AXIS_TKEEP,
    SLOT_6_AXIS_TLAST,
    SLOT_6_AXIS_TID,
    SLOT_6_AXIS_TDEST,
    SLOT_6_AXIS_TUSER,
    SLOT_7_AXI_ACLK,
    SLOT_7_AXI_ARESETN,
    SLOT_7_AXI_AWID,
    SLOT_7_AXI_AWADDR,
    SLOT_7_AXI_AWLEN,
    SLOT_7_AXI_AWPROT,
    SLOT_7_AXI_AWSIZE,
    SLOT_7_AXI_AWBURST,
    SLOT_7_AXI_AWCACHE,
    SLOT_7_AXI_AWLOCK,
    SLOT_7_AXI_AWVALID,
    SLOT_7_AXI_AWREADY,
    SLOT_7_AXI_WDATA,
    SLOT_7_AXI_WSTRB,
    SLOT_7_AXI_WLAST,
    SLOT_7_AXI_WVALID,
    SLOT_7_AXI_WREADY,
    SLOT_7_AXI_BID,
    SLOT_7_AXI_BRESP,
    SLOT_7_AXI_BVALID,
    SLOT_7_AXI_BREADY,
    SLOT_7_AXI_ARID,
    SLOT_7_AXI_ARADDR,
    SLOT_7_AXI_ARLEN,
    SLOT_7_AXI_ARSIZE,
    SLOT_7_AXI_ARBURST,
    SLOT_7_AXI_ARPROT,
    SLOT_7_AXI_ARCACHE,
    SLOT_7_AXI_ARLOCK,
    SLOT_7_AXI_ARVALID,
    SLOT_7_AXI_ARREADY,
    SLOT_7_AXI_RID,
    SLOT_7_AXI_RDATA,
    SLOT_7_AXI_RRESP,
    SLOT_7_AXI_RLAST,
    SLOT_7_AXI_RVALID,
    SLOT_7_AXI_RREADY,
    SLOT_7_AXIS_ACLK,
    SLOT_7_AXIS_ARESETN,
    SLOT_7_AXIS_TVALID,
    SLOT_7_AXIS_TREADY,
    SLOT_7_AXIS_TDATA,
    SLOT_7_AXIS_TSTRB,
    SLOT_7_AXIS_TKEEP,
    SLOT_7_AXIS_TLAST,
    SLOT_7_AXIS_TID,
    SLOT_7_AXIS_TDEST,
    SLOT_7_AXIS_TUSER,
    EXT_CLK_0,
    EXT_RSTN_0,
    EXT_EVENT_0_CNT_START,
    EXT_EVENT_0_CNT_STOP,
    EXT_EVENT_0,
    EXT_CLK_1,
    EXT_RSTN_1,
    EXT_EVENT_1_CNT_START,
    EXT_EVENT_1_CNT_STOP,
    EXT_EVENT_1,
    EXT_CLK_2,
    EXT_RSTN_2,
    EXT_EVENT_2_CNT_START,
    EXT_EVENT_2_CNT_STOP,
    EXT_EVENT_2,
    EXT_CLK_3,
    EXT_RSTN_3,
    EXT_EVENT_3_CNT_START,
    EXT_EVENT_3_CNT_STOP,
    EXT_EVENT_3,
    EXT_CLK_4,
    EXT_RSTN_4,
    EXT_EVENT_4_CNT_START,
    EXT_EVENT_4_CNT_STOP,
    EXT_EVENT_4,
    EXT_CLK_5,
    EXT_RSTN_5,
    EXT_EVENT_5_CNT_START,
    EXT_EVENT_5_CNT_STOP,
    EXT_EVENT_5,
    EXT_CLK_6,
    EXT_RSTN_6,
    EXT_EVENT_6_CNT_START,
    EXT_EVENT_6_CNT_STOP,
    EXT_EVENT_6,
    EXT_CLK_7,
    EXT_RSTN_7,
    EXT_EVENT_7_CNT_START,
    EXT_EVENT_7_CNT_STOP,
    EXT_EVENT_7,
    SLOT_0_EXT_TRIG,
    SLOT_1_EXT_TRIG,
    SLOT_2_EXT_TRIG,
    SLOT_3_EXT_TRIG,
    SLOT_4_EXT_TRIG,
    SLOT_5_EXT_TRIG,
    SLOT_6_EXT_TRIG,
    SLOT_7_EXT_TRIG,
    CAPTURE_EVENT,
    RESET_EVENT,
    M_AXIS_ACLK,
    M_AXIS_ARESETN,
    M_AXIS_TDATA,
    M_AXIS_TSTRB,
    M_AXIS_TVALID,
    M_AXIS_TID,
    M_AXIS_TREADY,
    CORE_ACLK,
    CORE_ARESETN,
    INTERRUPT
  );
  input S_AXI_ACLK;
  input S_AXI_ARESETN;
  input [15:0] S_AXI_AWADDR;
  input S_AXI_AWVALID;
  output S_AXI_AWREADY;
  input [31:0] S_AXI_WDATA;
  input [3:0] S_AXI_WSTRB;
  input S_AXI_WVALID;
  output S_AXI_WREADY;
  output [1:0] S_AXI_BRESP;
  output S_AXI_BVALID;
  input S_AXI_BREADY;
  input [15:0] S_AXI_ARADDR;
  input S_AXI_ARVALID;
  output S_AXI_ARREADY;
  output [31:0] S_AXI_RDATA;
  output [1:0] S_AXI_RRESP;
  output S_AXI_RVALID;
  input S_AXI_RREADY;
  input SLOT_0_AXI_ACLK;
  input SLOT_0_AXI_ARESETN;
  input [0:0] SLOT_0_AXI_AWID;
  input [31:0] SLOT_0_AXI_AWADDR;
  input [7:0] SLOT_0_AXI_AWLEN;
  input [2:0] SLOT_0_AXI_AWPROT;
  input [2:0] SLOT_0_AXI_AWSIZE;
  input [1:0] SLOT_0_AXI_AWBURST;
  input [3:0] SLOT_0_AXI_AWCACHE;
  input SLOT_0_AXI_AWLOCK;
  input SLOT_0_AXI_AWVALID;
  input SLOT_0_AXI_AWREADY;
  input [63:0] SLOT_0_AXI_WDATA;
  input [7:0] SLOT_0_AXI_WSTRB;
  input SLOT_0_AXI_WLAST;
  input SLOT_0_AXI_WVALID;
  input SLOT_0_AXI_WREADY;
  input [0:0] SLOT_0_AXI_BID;
  input [1:0] SLOT_0_AXI_BRESP;
  input SLOT_0_AXI_BVALID;
  input SLOT_0_AXI_BREADY;
  input [0:0] SLOT_0_AXI_ARID;
  input [31:0] SLOT_0_AXI_ARADDR;
  input [7:0] SLOT_0_AXI_ARLEN;
  input [2:0] SLOT_0_AXI_ARSIZE;
  input [1:0] SLOT_0_AXI_ARBURST;
  input [2:0] SLOT_0_AXI_ARPROT;
  input [3:0] SLOT_0_AXI_ARCACHE;
  input SLOT_0_AXI_ARLOCK;
  input SLOT_0_AXI_ARVALID;
  input SLOT_0_AXI_ARREADY;
  input [0:0] SLOT_0_AXI_RID;
  input [63:0] SLOT_0_AXI_RDATA;
  input [1:0] SLOT_0_AXI_RRESP;
  input SLOT_0_AXI_RLAST;
  input SLOT_0_AXI_RVALID;
  input SLOT_0_AXI_RREADY;
  input SLOT_0_AXIS_ACLK;
  input SLOT_0_AXIS_ARESETN;
  input SLOT_0_AXIS_TVALID;
  input SLOT_0_AXIS_TREADY;
  input [31:0] SLOT_0_AXIS_TDATA;
  input [3:0] SLOT_0_AXIS_TSTRB;
  input [3:0] SLOT_0_AXIS_TKEEP;
  input SLOT_0_AXIS_TLAST;
  input [0:0] SLOT_0_AXIS_TID;
  input [0:0] SLOT_0_AXIS_TDEST;
  input [0:0] SLOT_0_AXIS_TUSER;
  input SLOT_1_AXI_ACLK;
  input SLOT_1_AXI_ARESETN;
  input [0:0] SLOT_1_AXI_AWID;
  input [31:0] SLOT_1_AXI_AWADDR;
  input [7:0] SLOT_1_AXI_AWLEN;
  input [2:0] SLOT_1_AXI_AWPROT;
  input [2:0] SLOT_1_AXI_AWSIZE;
  input [1:0] SLOT_1_AXI_AWBURST;
  input [3:0] SLOT_1_AXI_AWCACHE;
  input SLOT_1_AXI_AWLOCK;
  input SLOT_1_AXI_AWVALID;
  input SLOT_1_AXI_AWREADY;
  input [31:0] SLOT_1_AXI_WDATA;
  input [3:0] SLOT_1_AXI_WSTRB;
  input SLOT_1_AXI_WLAST;
  input SLOT_1_AXI_WVALID;
  input SLOT_1_AXI_WREADY;
  input [0:0] SLOT_1_AXI_BID;
  input [1:0] SLOT_1_AXI_BRESP;
  input SLOT_1_AXI_BVALID;
  input SLOT_1_AXI_BREADY;
  input [0:0] SLOT_1_AXI_ARID;
  input [31:0] SLOT_1_AXI_ARADDR;
  input [7:0] SLOT_1_AXI_ARLEN;
  input [2:0] SLOT_1_AXI_ARSIZE;
  input [1:0] SLOT_1_AXI_ARBURST;
  input [2:0] SLOT_1_AXI_ARPROT;
  input [3:0] SLOT_1_AXI_ARCACHE;
  input SLOT_1_AXI_ARLOCK;
  input SLOT_1_AXI_ARVALID;
  input SLOT_1_AXI_ARREADY;
  input [0:0] SLOT_1_AXI_RID;
  input [31:0] SLOT_1_AXI_RDATA;
  input [1:0] SLOT_1_AXI_RRESP;
  input SLOT_1_AXI_RLAST;
  input SLOT_1_AXI_RVALID;
  input SLOT_1_AXI_RREADY;
  input SLOT_1_AXIS_ACLK;
  input SLOT_1_AXIS_ARESETN;
  input SLOT_1_AXIS_TVALID;
  input SLOT_1_AXIS_TREADY;
  input [31:0] SLOT_1_AXIS_TDATA;
  input [3:0] SLOT_1_AXIS_TSTRB;
  input [3:0] SLOT_1_AXIS_TKEEP;
  input SLOT_1_AXIS_TLAST;
  input [0:0] SLOT_1_AXIS_TID;
  input [0:0] SLOT_1_AXIS_TDEST;
  input [0:0] SLOT_1_AXIS_TUSER;
  input SLOT_2_AXI_ACLK;
  input SLOT_2_AXI_ARESETN;
  input [0:0] SLOT_2_AXI_AWID;
  input [31:0] SLOT_2_AXI_AWADDR;
  input [7:0] SLOT_2_AXI_AWLEN;
  input [2:0] SLOT_2_AXI_AWPROT;
  input [2:0] SLOT_2_AXI_AWSIZE;
  input [1:0] SLOT_2_AXI_AWBURST;
  input [3:0] SLOT_2_AXI_AWCACHE;
  input SLOT_2_AXI_AWLOCK;
  input SLOT_2_AXI_AWVALID;
  input SLOT_2_AXI_AWREADY;
  input [31:0] SLOT_2_AXI_WDATA;
  input [3:0] SLOT_2_AXI_WSTRB;
  input SLOT_2_AXI_WLAST;
  input SLOT_2_AXI_WVALID;
  input SLOT_2_AXI_WREADY;
  input [0:0] SLOT_2_AXI_BID;
  input [1:0] SLOT_2_AXI_BRESP;
  input SLOT_2_AXI_BVALID;
  input SLOT_2_AXI_BREADY;
  input [0:0] SLOT_2_AXI_ARID;
  input [31:0] SLOT_2_AXI_ARADDR;
  input [7:0] SLOT_2_AXI_ARLEN;
  input [2:0] SLOT_2_AXI_ARSIZE;
  input [1:0] SLOT_2_AXI_ARBURST;
  input [2:0] SLOT_2_AXI_ARPROT;
  input [3:0] SLOT_2_AXI_ARCACHE;
  input SLOT_2_AXI_ARLOCK;
  input SLOT_2_AXI_ARVALID;
  input SLOT_2_AXI_ARREADY;
  input [0:0] SLOT_2_AXI_RID;
  input [31:0] SLOT_2_AXI_RDATA;
  input [1:0] SLOT_2_AXI_RRESP;
  input SLOT_2_AXI_RLAST;
  input SLOT_2_AXI_RVALID;
  input SLOT_2_AXI_RREADY;
  input SLOT_2_AXIS_ACLK;
  input SLOT_2_AXIS_ARESETN;
  input SLOT_2_AXIS_TVALID;
  input SLOT_2_AXIS_TREADY;
  input [31:0] SLOT_2_AXIS_TDATA;
  input [3:0] SLOT_2_AXIS_TSTRB;
  input [3:0] SLOT_2_AXIS_TKEEP;
  input SLOT_2_AXIS_TLAST;
  input [0:0] SLOT_2_AXIS_TID;
  input [0:0] SLOT_2_AXIS_TDEST;
  input [0:0] SLOT_2_AXIS_TUSER;
  input SLOT_3_AXI_ACLK;
  input SLOT_3_AXI_ARESETN;
  input [0:0] SLOT_3_AXI_AWID;
  input [31:0] SLOT_3_AXI_AWADDR;
  input [7:0] SLOT_3_AXI_AWLEN;
  input [2:0] SLOT_3_AXI_AWPROT;
  input [2:0] SLOT_3_AXI_AWSIZE;
  input [1:0] SLOT_3_AXI_AWBURST;
  input [3:0] SLOT_3_AXI_AWCACHE;
  input SLOT_3_AXI_AWLOCK;
  input SLOT_3_AXI_AWVALID;
  input SLOT_3_AXI_AWREADY;
  input [31:0] SLOT_3_AXI_WDATA;
  input [3:0] SLOT_3_AXI_WSTRB;
  input SLOT_3_AXI_WLAST;
  input SLOT_3_AXI_WVALID;
  input SLOT_3_AXI_WREADY;
  input [0:0] SLOT_3_AXI_BID;
  input [1:0] SLOT_3_AXI_BRESP;
  input SLOT_3_AXI_BVALID;
  input SLOT_3_AXI_BREADY;
  input [0:0] SLOT_3_AXI_ARID;
  input [31:0] SLOT_3_AXI_ARADDR;
  input [7:0] SLOT_3_AXI_ARLEN;
  input [2:0] SLOT_3_AXI_ARSIZE;
  input [1:0] SLOT_3_AXI_ARBURST;
  input [2:0] SLOT_3_AXI_ARPROT;
  input [3:0] SLOT_3_AXI_ARCACHE;
  input SLOT_3_AXI_ARLOCK;
  input SLOT_3_AXI_ARVALID;
  input SLOT_3_AXI_ARREADY;
  input [0:0] SLOT_3_AXI_RID;
  input [31:0] SLOT_3_AXI_RDATA;
  input [1:0] SLOT_3_AXI_RRESP;
  input SLOT_3_AXI_RLAST;
  input SLOT_3_AXI_RVALID;
  input SLOT_3_AXI_RREADY;
  input SLOT_3_AXIS_ACLK;
  input SLOT_3_AXIS_ARESETN;
  input SLOT_3_AXIS_TVALID;
  input SLOT_3_AXIS_TREADY;
  input [31:0] SLOT_3_AXIS_TDATA;
  input [3:0] SLOT_3_AXIS_TSTRB;
  input [3:0] SLOT_3_AXIS_TKEEP;
  input SLOT_3_AXIS_TLAST;
  input [0:0] SLOT_3_AXIS_TID;
  input [0:0] SLOT_3_AXIS_TDEST;
  input [0:0] SLOT_3_AXIS_TUSER;
  input SLOT_4_AXI_ACLK;
  input SLOT_4_AXI_ARESETN;
  input [0:0] SLOT_4_AXI_AWID;
  input [31:0] SLOT_4_AXI_AWADDR;
  input [7:0] SLOT_4_AXI_AWLEN;
  input [2:0] SLOT_4_AXI_AWPROT;
  input [2:0] SLOT_4_AXI_AWSIZE;
  input [1:0] SLOT_4_AXI_AWBURST;
  input [3:0] SLOT_4_AXI_AWCACHE;
  input SLOT_4_AXI_AWLOCK;
  input SLOT_4_AXI_AWVALID;
  input SLOT_4_AXI_AWREADY;
  input [31:0] SLOT_4_AXI_WDATA;
  input [3:0] SLOT_4_AXI_WSTRB;
  input SLOT_4_AXI_WLAST;
  input SLOT_4_AXI_WVALID;
  input SLOT_4_AXI_WREADY;
  input [0:0] SLOT_4_AXI_BID;
  input [1:0] SLOT_4_AXI_BRESP;
  input SLOT_4_AXI_BVALID;
  input SLOT_4_AXI_BREADY;
  input [0:0] SLOT_4_AXI_ARID;
  input [31:0] SLOT_4_AXI_ARADDR;
  input [7:0] SLOT_4_AXI_ARLEN;
  input [2:0] SLOT_4_AXI_ARSIZE;
  input [1:0] SLOT_4_AXI_ARBURST;
  input [2:0] SLOT_4_AXI_ARPROT;
  input [3:0] SLOT_4_AXI_ARCACHE;
  input SLOT_4_AXI_ARLOCK;
  input SLOT_4_AXI_ARVALID;
  input SLOT_4_AXI_ARREADY;
  input [0:0] SLOT_4_AXI_RID;
  input [31:0] SLOT_4_AXI_RDATA;
  input [1:0] SLOT_4_AXI_RRESP;
  input SLOT_4_AXI_RLAST;
  input SLOT_4_AXI_RVALID;
  input SLOT_4_AXI_RREADY;
  input SLOT_4_AXIS_ACLK;
  input SLOT_4_AXIS_ARESETN;
  input SLOT_4_AXIS_TVALID;
  input SLOT_4_AXIS_TREADY;
  input [31:0] SLOT_4_AXIS_TDATA;
  input [3:0] SLOT_4_AXIS_TSTRB;
  input [3:0] SLOT_4_AXIS_TKEEP;
  input SLOT_4_AXIS_TLAST;
  input [0:0] SLOT_4_AXIS_TID;
  input [0:0] SLOT_4_AXIS_TDEST;
  input [0:0] SLOT_4_AXIS_TUSER;
  input SLOT_5_AXI_ACLK;
  input SLOT_5_AXI_ARESETN;
  input [0:0] SLOT_5_AXI_AWID;
  input [31:0] SLOT_5_AXI_AWADDR;
  input [7:0] SLOT_5_AXI_AWLEN;
  input [2:0] SLOT_5_AXI_AWPROT;
  input [2:0] SLOT_5_AXI_AWSIZE;
  input [1:0] SLOT_5_AXI_AWBURST;
  input [3:0] SLOT_5_AXI_AWCACHE;
  input SLOT_5_AXI_AWLOCK;
  input SLOT_5_AXI_AWVALID;
  input SLOT_5_AXI_AWREADY;
  input [31:0] SLOT_5_AXI_WDATA;
  input [3:0] SLOT_5_AXI_WSTRB;
  input SLOT_5_AXI_WLAST;
  input SLOT_5_AXI_WVALID;
  input SLOT_5_AXI_WREADY;
  input [0:0] SLOT_5_AXI_BID;
  input [1:0] SLOT_5_AXI_BRESP;
  input SLOT_5_AXI_BVALID;
  input SLOT_5_AXI_BREADY;
  input [0:0] SLOT_5_AXI_ARID;
  input [31:0] SLOT_5_AXI_ARADDR;
  input [7:0] SLOT_5_AXI_ARLEN;
  input [2:0] SLOT_5_AXI_ARSIZE;
  input [1:0] SLOT_5_AXI_ARBURST;
  input [2:0] SLOT_5_AXI_ARPROT;
  input [3:0] SLOT_5_AXI_ARCACHE;
  input SLOT_5_AXI_ARLOCK;
  input SLOT_5_AXI_ARVALID;
  input SLOT_5_AXI_ARREADY;
  input [0:0] SLOT_5_AXI_RID;
  input [31:0] SLOT_5_AXI_RDATA;
  input [1:0] SLOT_5_AXI_RRESP;
  input SLOT_5_AXI_RLAST;
  input SLOT_5_AXI_RVALID;
  input SLOT_5_AXI_RREADY;
  input SLOT_5_AXIS_ACLK;
  input SLOT_5_AXIS_ARESETN;
  input SLOT_5_AXIS_TVALID;
  input SLOT_5_AXIS_TREADY;
  input [31:0] SLOT_5_AXIS_TDATA;
  input [3:0] SLOT_5_AXIS_TSTRB;
  input [3:0] SLOT_5_AXIS_TKEEP;
  input SLOT_5_AXIS_TLAST;
  input [0:0] SLOT_5_AXIS_TID;
  input [0:0] SLOT_5_AXIS_TDEST;
  input [0:0] SLOT_5_AXIS_TUSER;
  input SLOT_6_AXI_ACLK;
  input SLOT_6_AXI_ARESETN;
  input [0:0] SLOT_6_AXI_AWID;
  input [31:0] SLOT_6_AXI_AWADDR;
  input [7:0] SLOT_6_AXI_AWLEN;
  input [2:0] SLOT_6_AXI_AWPROT;
  input [2:0] SLOT_6_AXI_AWSIZE;
  input [1:0] SLOT_6_AXI_AWBURST;
  input [3:0] SLOT_6_AXI_AWCACHE;
  input SLOT_6_AXI_AWLOCK;
  input SLOT_6_AXI_AWVALID;
  input SLOT_6_AXI_AWREADY;
  input [31:0] SLOT_6_AXI_WDATA;
  input [3:0] SLOT_6_AXI_WSTRB;
  input SLOT_6_AXI_WLAST;
  input SLOT_6_AXI_WVALID;
  input SLOT_6_AXI_WREADY;
  input [0:0] SLOT_6_AXI_BID;
  input [1:0] SLOT_6_AXI_BRESP;
  input SLOT_6_AXI_BVALID;
  input SLOT_6_AXI_BREADY;
  input [0:0] SLOT_6_AXI_ARID;
  input [31:0] SLOT_6_AXI_ARADDR;
  input [7:0] SLOT_6_AXI_ARLEN;
  input [2:0] SLOT_6_AXI_ARSIZE;
  input [1:0] SLOT_6_AXI_ARBURST;
  input [2:0] SLOT_6_AXI_ARPROT;
  input [3:0] SLOT_6_AXI_ARCACHE;
  input SLOT_6_AXI_ARLOCK;
  input SLOT_6_AXI_ARVALID;
  input SLOT_6_AXI_ARREADY;
  input [0:0] SLOT_6_AXI_RID;
  input [31:0] SLOT_6_AXI_RDATA;
  input [1:0] SLOT_6_AXI_RRESP;
  input SLOT_6_AXI_RLAST;
  input SLOT_6_AXI_RVALID;
  input SLOT_6_AXI_RREADY;
  input SLOT_6_AXIS_ACLK;
  input SLOT_6_AXIS_ARESETN;
  input SLOT_6_AXIS_TVALID;
  input SLOT_6_AXIS_TREADY;
  input [31:0] SLOT_6_AXIS_TDATA;
  input [3:0] SLOT_6_AXIS_TSTRB;
  input [3:0] SLOT_6_AXIS_TKEEP;
  input SLOT_6_AXIS_TLAST;
  input [0:0] SLOT_6_AXIS_TID;
  input [0:0] SLOT_6_AXIS_TDEST;
  input [0:0] SLOT_6_AXIS_TUSER;
  input SLOT_7_AXI_ACLK;
  input SLOT_7_AXI_ARESETN;
  input [0:0] SLOT_7_AXI_AWID;
  input [31:0] SLOT_7_AXI_AWADDR;
  input [7:0] SLOT_7_AXI_AWLEN;
  input [2:0] SLOT_7_AXI_AWPROT;
  input [2:0] SLOT_7_AXI_AWSIZE;
  input [1:0] SLOT_7_AXI_AWBURST;
  input [3:0] SLOT_7_AXI_AWCACHE;
  input SLOT_7_AXI_AWLOCK;
  input SLOT_7_AXI_AWVALID;
  input SLOT_7_AXI_AWREADY;
  input [31:0] SLOT_7_AXI_WDATA;
  input [3:0] SLOT_7_AXI_WSTRB;
  input SLOT_7_AXI_WLAST;
  input SLOT_7_AXI_WVALID;
  input SLOT_7_AXI_WREADY;
  input [0:0] SLOT_7_AXI_BID;
  input [1:0] SLOT_7_AXI_BRESP;
  input SLOT_7_AXI_BVALID;
  input SLOT_7_AXI_BREADY;
  input [0:0] SLOT_7_AXI_ARID;
  input [31:0] SLOT_7_AXI_ARADDR;
  input [7:0] SLOT_7_AXI_ARLEN;
  input [2:0] SLOT_7_AXI_ARSIZE;
  input [1:0] SLOT_7_AXI_ARBURST;
  input [2:0] SLOT_7_AXI_ARPROT;
  input [3:0] SLOT_7_AXI_ARCACHE;
  input SLOT_7_AXI_ARLOCK;
  input SLOT_7_AXI_ARVALID;
  input SLOT_7_AXI_ARREADY;
  input [0:0] SLOT_7_AXI_RID;
  input [31:0] SLOT_7_AXI_RDATA;
  input [1:0] SLOT_7_AXI_RRESP;
  input SLOT_7_AXI_RLAST;
  input SLOT_7_AXI_RVALID;
  input SLOT_7_AXI_RREADY;
  input SLOT_7_AXIS_ACLK;
  input SLOT_7_AXIS_ARESETN;
  input SLOT_7_AXIS_TVALID;
  input SLOT_7_AXIS_TREADY;
  input [31:0] SLOT_7_AXIS_TDATA;
  input [3:0] SLOT_7_AXIS_TSTRB;
  input [3:0] SLOT_7_AXIS_TKEEP;
  input SLOT_7_AXIS_TLAST;
  input [0:0] SLOT_7_AXIS_TID;
  input [0:0] SLOT_7_AXIS_TDEST;
  input [0:0] SLOT_7_AXIS_TUSER;
  input EXT_CLK_0;
  input EXT_RSTN_0;
  input EXT_EVENT_0_CNT_START;
  input EXT_EVENT_0_CNT_STOP;
  input EXT_EVENT_0;
  input EXT_CLK_1;
  input EXT_RSTN_1;
  input EXT_EVENT_1_CNT_START;
  input EXT_EVENT_1_CNT_STOP;
  input EXT_EVENT_1;
  input EXT_CLK_2;
  input EXT_RSTN_2;
  input EXT_EVENT_2_CNT_START;
  input EXT_EVENT_2_CNT_STOP;
  input EXT_EVENT_2;
  input EXT_CLK_3;
  input EXT_RSTN_3;
  input EXT_EVENT_3_CNT_START;
  input EXT_EVENT_3_CNT_STOP;
  input EXT_EVENT_3;
  input EXT_CLK_4;
  input EXT_RSTN_4;
  input EXT_EVENT_4_CNT_START;
  input EXT_EVENT_4_CNT_STOP;
  input EXT_EVENT_4;
  input EXT_CLK_5;
  input EXT_RSTN_5;
  input EXT_EVENT_5_CNT_START;
  input EXT_EVENT_5_CNT_STOP;
  input EXT_EVENT_5;
  input EXT_CLK_6;
  input EXT_RSTN_6;
  input EXT_EVENT_6_CNT_START;
  input EXT_EVENT_6_CNT_STOP;
  input EXT_EVENT_6;
  input EXT_CLK_7;
  input EXT_RSTN_7;
  input EXT_EVENT_7_CNT_START;
  input EXT_EVENT_7_CNT_STOP;
  input EXT_EVENT_7;
  input SLOT_0_EXT_TRIG;
  input SLOT_1_EXT_TRIG;
  input SLOT_2_EXT_TRIG;
  input SLOT_3_EXT_TRIG;
  input SLOT_4_EXT_TRIG;
  input SLOT_5_EXT_TRIG;
  input SLOT_6_EXT_TRIG;
  input SLOT_7_EXT_TRIG;
  input CAPTURE_EVENT;
  input RESET_EVENT;
  input M_AXIS_ACLK;
  input M_AXIS_ARESETN;
  output [55:0] M_AXIS_TDATA;
  output [6:0] M_AXIS_TSTRB;
  output M_AXIS_TVALID;
  output [0:0] M_AXIS_TID;
  input M_AXIS_TREADY;
  input CORE_ACLK;
  input CORE_ARESETN;
  output INTERRUPT;

  axi_perf_mon
    #(
      .C_FAMILY ( "zynq" ),
      .C_INSTANCE ( "axi_perf_mon_0" ),
      .C_S_AXI_ADDR_WIDTH ( 16 ),
      .C_S_AXI_DATA_WIDTH ( 32 ),
      .C_NUM_MONITOR_SLOTS ( 1 ),
      .C_ENABLE_EVENT_COUNT ( 1 ),
      .C_NUM_OF_COUNTERS ( 4 ),
      .C_METRIC_COUNT_WIDTH ( 32 ),
      .C_GLOBAL_COUNT_WIDTH ( 64 ),
      .C_METRICS_SAMPLE_COUNT_WIDTH ( 64 ),
      .C_MAX_OUTSTAND_DEPTH ( 1 ),
      .C_MAX_REORDER_DEPTH ( 1 ),
      .C_SLOT_0_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_0_AXI_DATA_WIDTH ( 64 ),
      .C_SLOT_0_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_0_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_0_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_0_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_0_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_0_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_0_FIFO_ENABLE ( 1 ),
      .C_SLOT_1_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_1_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_1_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_1_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_1_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_1_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_1_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_1_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_1_FIFO_ENABLE ( 1 ),
      .C_SLOT_2_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_2_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_2_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_2_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_2_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_2_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_2_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_2_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_2_FIFO_ENABLE ( 1 ),
      .C_SLOT_3_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_3_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_3_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_3_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_3_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_3_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_3_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_3_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_3_FIFO_ENABLE ( 1 ),
      .C_SLOT_4_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_4_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_4_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_4_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_4_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_4_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_4_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_4_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_4_FIFO_ENABLE ( 1 ),
      .C_SLOT_5_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_5_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_5_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_5_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_5_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_5_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_5_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_5_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_5_FIFO_ENABLE ( 1 ),
      .C_SLOT_6_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_6_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_6_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_6_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_6_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_6_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_6_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_6_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_6_FIFO_ENABLE ( 1 ),
      .C_SLOT_7_AXI_ADDR_WIDTH ( 32 ),
      .C_SLOT_7_AXI_DATA_WIDTH ( 32 ),
      .C_SLOT_7_AXI_ID_WIDTH ( 1 ),
      .C_SLOT_7_AXI_PROTOCOL ( "AXI4MM" ),
      .C_SLOT_7_AXIS_TDATA_WIDTH ( 32 ),
      .C_SLOT_7_AXIS_TID_WIDTH ( 1 ),
      .C_SLOT_7_AXIS_TDEST_WIDTH ( 1 ),
      .C_SLOT_7_AXIS_TUSER_WIDTH ( 1 ),
      .C_SLOT_7_FIFO_ENABLE ( 1 ),
      .C_REG_ALL_MONITOR_SIGNALS ( 0 ),
      .C_EXT_EVENT0_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT1_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT2_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT3_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT4_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT5_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT6_FIFO_ENABLE ( 1 ),
      .C_EXT_EVENT7_FIFO_ENABLE ( 1 ),
      .C_ENABLE_EVENT_LOG ( 0 ),
      .C_FIFO_AXIS_DEPTH ( 32 ),
      .C_FIFO_AXIS_TDATA_WIDTH ( 56 ),
      .C_FIFO_AXIS_TID_WIDTH ( 1 ),
      .C_AXI4LITE_CORE_CLK_ASYNC ( 1 ),
      .C_HAVE_SAMPLED_METRIC_CNT ( 0 ),
      .C_FIFO_AXIS_SYNC ( 0 ),
      .C_SHOW_AXI_IDS ( 0 ),
      .C_SHOW_AXI_LEN ( 0 ),
      .C_SHOW_AXIS_TID ( 0 ),
      .C_SHOW_AXIS_TDEST ( 0 ),
      .C_SHOW_AXIS_TUSER ( 0 )
    )
    axi_perf_mon_0 (
      .S_AXI_ACLK ( S_AXI_ACLK ),
      .S_AXI_ARESETN ( S_AXI_ARESETN ),
      .S_AXI_AWADDR ( S_AXI_AWADDR ),
      .S_AXI_AWVALID ( S_AXI_AWVALID ),
      .S_AXI_AWREADY ( S_AXI_AWREADY ),
      .S_AXI_WDATA ( S_AXI_WDATA ),
      .S_AXI_WSTRB ( S_AXI_WSTRB ),
      .S_AXI_WVALID ( S_AXI_WVALID ),
      .S_AXI_WREADY ( S_AXI_WREADY ),
      .S_AXI_BRESP ( S_AXI_BRESP ),
      .S_AXI_BVALID ( S_AXI_BVALID ),
      .S_AXI_BREADY ( S_AXI_BREADY ),
      .S_AXI_ARADDR ( S_AXI_ARADDR ),
      .S_AXI_ARVALID ( S_AXI_ARVALID ),
      .S_AXI_ARREADY ( S_AXI_ARREADY ),
      .S_AXI_RDATA ( S_AXI_RDATA ),
      .S_AXI_RRESP ( S_AXI_RRESP ),
      .S_AXI_RVALID ( S_AXI_RVALID ),
      .S_AXI_RREADY ( S_AXI_RREADY ),
      .SLOT_0_AXI_ACLK ( SLOT_0_AXI_ACLK ),
      .SLOT_0_AXI_ARESETN ( SLOT_0_AXI_ARESETN ),
      .SLOT_0_AXI_AWID ( SLOT_0_AXI_AWID ),
      .SLOT_0_AXI_AWADDR ( SLOT_0_AXI_AWADDR ),
      .SLOT_0_AXI_AWLEN ( SLOT_0_AXI_AWLEN ),
      .SLOT_0_AXI_AWPROT ( SLOT_0_AXI_AWPROT ),
      .SLOT_0_AXI_AWSIZE ( SLOT_0_AXI_AWSIZE ),
      .SLOT_0_AXI_AWBURST ( SLOT_0_AXI_AWBURST ),
      .SLOT_0_AXI_AWCACHE ( SLOT_0_AXI_AWCACHE ),
      .SLOT_0_AXI_AWLOCK ( SLOT_0_AXI_AWLOCK ),
      .SLOT_0_AXI_AWVALID ( SLOT_0_AXI_AWVALID ),
      .SLOT_0_AXI_AWREADY ( SLOT_0_AXI_AWREADY ),
      .SLOT_0_AXI_WDATA ( SLOT_0_AXI_WDATA ),
      .SLOT_0_AXI_WSTRB ( SLOT_0_AXI_WSTRB ),
      .SLOT_0_AXI_WLAST ( SLOT_0_AXI_WLAST ),
      .SLOT_0_AXI_WVALID ( SLOT_0_AXI_WVALID ),
      .SLOT_0_AXI_WREADY ( SLOT_0_AXI_WREADY ),
      .SLOT_0_AXI_BID ( SLOT_0_AXI_BID ),
      .SLOT_0_AXI_BRESP ( SLOT_0_AXI_BRESP ),
      .SLOT_0_AXI_BVALID ( SLOT_0_AXI_BVALID ),
      .SLOT_0_AXI_BREADY ( SLOT_0_AXI_BREADY ),
      .SLOT_0_AXI_ARID ( SLOT_0_AXI_ARID ),
      .SLOT_0_AXI_ARADDR ( SLOT_0_AXI_ARADDR ),
      .SLOT_0_AXI_ARLEN ( SLOT_0_AXI_ARLEN ),
      .SLOT_0_AXI_ARSIZE ( SLOT_0_AXI_ARSIZE ),
      .SLOT_0_AXI_ARBURST ( SLOT_0_AXI_ARBURST ),
      .SLOT_0_AXI_ARPROT ( SLOT_0_AXI_ARPROT ),
      .SLOT_0_AXI_ARCACHE ( SLOT_0_AXI_ARCACHE ),
      .SLOT_0_AXI_ARLOCK ( SLOT_0_AXI_ARLOCK ),
      .SLOT_0_AXI_ARVALID ( SLOT_0_AXI_ARVALID ),
      .SLOT_0_AXI_ARREADY ( SLOT_0_AXI_ARREADY ),
      .SLOT_0_AXI_RID ( SLOT_0_AXI_RID ),
      .SLOT_0_AXI_RDATA ( SLOT_0_AXI_RDATA ),
      .SLOT_0_AXI_RRESP ( SLOT_0_AXI_RRESP ),
      .SLOT_0_AXI_RLAST ( SLOT_0_AXI_RLAST ),
      .SLOT_0_AXI_RVALID ( SLOT_0_AXI_RVALID ),
      .SLOT_0_AXI_RREADY ( SLOT_0_AXI_RREADY ),
      .SLOT_0_AXIS_ACLK ( SLOT_0_AXIS_ACLK ),
      .SLOT_0_AXIS_ARESETN ( SLOT_0_AXIS_ARESETN ),
      .SLOT_0_AXIS_TVALID ( SLOT_0_AXIS_TVALID ),
      .SLOT_0_AXIS_TREADY ( SLOT_0_AXIS_TREADY ),
      .SLOT_0_AXIS_TDATA ( SLOT_0_AXIS_TDATA ),
      .SLOT_0_AXIS_TSTRB ( SLOT_0_AXIS_TSTRB ),
      .SLOT_0_AXIS_TKEEP ( SLOT_0_AXIS_TKEEP ),
      .SLOT_0_AXIS_TLAST ( SLOT_0_AXIS_TLAST ),
      .SLOT_0_AXIS_TID ( SLOT_0_AXIS_TID ),
      .SLOT_0_AXIS_TDEST ( SLOT_0_AXIS_TDEST ),
      .SLOT_0_AXIS_TUSER ( SLOT_0_AXIS_TUSER ),
      .SLOT_1_AXI_ACLK ( SLOT_1_AXI_ACLK ),
      .SLOT_1_AXI_ARESETN ( SLOT_1_AXI_ARESETN ),
      .SLOT_1_AXI_AWID ( SLOT_1_AXI_AWID ),
      .SLOT_1_AXI_AWADDR ( SLOT_1_AXI_AWADDR ),
      .SLOT_1_AXI_AWLEN ( SLOT_1_AXI_AWLEN ),
      .SLOT_1_AXI_AWPROT ( SLOT_1_AXI_AWPROT ),
      .SLOT_1_AXI_AWSIZE ( SLOT_1_AXI_AWSIZE ),
      .SLOT_1_AXI_AWBURST ( SLOT_1_AXI_AWBURST ),
      .SLOT_1_AXI_AWCACHE ( SLOT_1_AXI_AWCACHE ),
      .SLOT_1_AXI_AWLOCK ( SLOT_1_AXI_AWLOCK ),
      .SLOT_1_AXI_AWVALID ( SLOT_1_AXI_AWVALID ),
      .SLOT_1_AXI_AWREADY ( SLOT_1_AXI_AWREADY ),
      .SLOT_1_AXI_WDATA ( SLOT_1_AXI_WDATA ),
      .SLOT_1_AXI_WSTRB ( SLOT_1_AXI_WSTRB ),
      .SLOT_1_AXI_WLAST ( SLOT_1_AXI_WLAST ),
      .SLOT_1_AXI_WVALID ( SLOT_1_AXI_WVALID ),
      .SLOT_1_AXI_WREADY ( SLOT_1_AXI_WREADY ),
      .SLOT_1_AXI_BID ( SLOT_1_AXI_BID ),
      .SLOT_1_AXI_BRESP ( SLOT_1_AXI_BRESP ),
      .SLOT_1_AXI_BVALID ( SLOT_1_AXI_BVALID ),
      .SLOT_1_AXI_BREADY ( SLOT_1_AXI_BREADY ),
      .SLOT_1_AXI_ARID ( SLOT_1_AXI_ARID ),
      .SLOT_1_AXI_ARADDR ( SLOT_1_AXI_ARADDR ),
      .SLOT_1_AXI_ARLEN ( SLOT_1_AXI_ARLEN ),
      .SLOT_1_AXI_ARSIZE ( SLOT_1_AXI_ARSIZE ),
      .SLOT_1_AXI_ARBURST ( SLOT_1_AXI_ARBURST ),
      .SLOT_1_AXI_ARPROT ( SLOT_1_AXI_ARPROT ),
      .SLOT_1_AXI_ARCACHE ( SLOT_1_AXI_ARCACHE ),
      .SLOT_1_AXI_ARLOCK ( SLOT_1_AXI_ARLOCK ),
      .SLOT_1_AXI_ARVALID ( SLOT_1_AXI_ARVALID ),
      .SLOT_1_AXI_ARREADY ( SLOT_1_AXI_ARREADY ),
      .SLOT_1_AXI_RID ( SLOT_1_AXI_RID ),
      .SLOT_1_AXI_RDATA ( SLOT_1_AXI_RDATA ),
      .SLOT_1_AXI_RRESP ( SLOT_1_AXI_RRESP ),
      .SLOT_1_AXI_RLAST ( SLOT_1_AXI_RLAST ),
      .SLOT_1_AXI_RVALID ( SLOT_1_AXI_RVALID ),
      .SLOT_1_AXI_RREADY ( SLOT_1_AXI_RREADY ),
      .SLOT_1_AXIS_ACLK ( SLOT_1_AXIS_ACLK ),
      .SLOT_1_AXIS_ARESETN ( SLOT_1_AXIS_ARESETN ),
      .SLOT_1_AXIS_TVALID ( SLOT_1_AXIS_TVALID ),
      .SLOT_1_AXIS_TREADY ( SLOT_1_AXIS_TREADY ),
      .SLOT_1_AXIS_TDATA ( SLOT_1_AXIS_TDATA ),
      .SLOT_1_AXIS_TSTRB ( SLOT_1_AXIS_TSTRB ),
      .SLOT_1_AXIS_TKEEP ( SLOT_1_AXIS_TKEEP ),
      .SLOT_1_AXIS_TLAST ( SLOT_1_AXIS_TLAST ),
      .SLOT_1_AXIS_TID ( SLOT_1_AXIS_TID ),
      .SLOT_1_AXIS_TDEST ( SLOT_1_AXIS_TDEST ),
      .SLOT_1_AXIS_TUSER ( SLOT_1_AXIS_TUSER ),
      .SLOT_2_AXI_ACLK ( SLOT_2_AXI_ACLK ),
      .SLOT_2_AXI_ARESETN ( SLOT_2_AXI_ARESETN ),
      .SLOT_2_AXI_AWID ( SLOT_2_AXI_AWID ),
      .SLOT_2_AXI_AWADDR ( SLOT_2_AXI_AWADDR ),
      .SLOT_2_AXI_AWLEN ( SLOT_2_AXI_AWLEN ),
      .SLOT_2_AXI_AWPROT ( SLOT_2_AXI_AWPROT ),
      .SLOT_2_AXI_AWSIZE ( SLOT_2_AXI_AWSIZE ),
      .SLOT_2_AXI_AWBURST ( SLOT_2_AXI_AWBURST ),
      .SLOT_2_AXI_AWCACHE ( SLOT_2_AXI_AWCACHE ),
      .SLOT_2_AXI_AWLOCK ( SLOT_2_AXI_AWLOCK ),
      .SLOT_2_AXI_AWVALID ( SLOT_2_AXI_AWVALID ),
      .SLOT_2_AXI_AWREADY ( SLOT_2_AXI_AWREADY ),
      .SLOT_2_AXI_WDATA ( SLOT_2_AXI_WDATA ),
      .SLOT_2_AXI_WSTRB ( SLOT_2_AXI_WSTRB ),
      .SLOT_2_AXI_WLAST ( SLOT_2_AXI_WLAST ),
      .SLOT_2_AXI_WVALID ( SLOT_2_AXI_WVALID ),
      .SLOT_2_AXI_WREADY ( SLOT_2_AXI_WREADY ),
      .SLOT_2_AXI_BID ( SLOT_2_AXI_BID ),
      .SLOT_2_AXI_BRESP ( SLOT_2_AXI_BRESP ),
      .SLOT_2_AXI_BVALID ( SLOT_2_AXI_BVALID ),
      .SLOT_2_AXI_BREADY ( SLOT_2_AXI_BREADY ),
      .SLOT_2_AXI_ARID ( SLOT_2_AXI_ARID ),
      .SLOT_2_AXI_ARADDR ( SLOT_2_AXI_ARADDR ),
      .SLOT_2_AXI_ARLEN ( SLOT_2_AXI_ARLEN ),
      .SLOT_2_AXI_ARSIZE ( SLOT_2_AXI_ARSIZE ),
      .SLOT_2_AXI_ARBURST ( SLOT_2_AXI_ARBURST ),
      .SLOT_2_AXI_ARPROT ( SLOT_2_AXI_ARPROT ),
      .SLOT_2_AXI_ARCACHE ( SLOT_2_AXI_ARCACHE ),
      .SLOT_2_AXI_ARLOCK ( SLOT_2_AXI_ARLOCK ),
      .SLOT_2_AXI_ARVALID ( SLOT_2_AXI_ARVALID ),
      .SLOT_2_AXI_ARREADY ( SLOT_2_AXI_ARREADY ),
      .SLOT_2_AXI_RID ( SLOT_2_AXI_RID ),
      .SLOT_2_AXI_RDATA ( SLOT_2_AXI_RDATA ),
      .SLOT_2_AXI_RRESP ( SLOT_2_AXI_RRESP ),
      .SLOT_2_AXI_RLAST ( SLOT_2_AXI_RLAST ),
      .SLOT_2_AXI_RVALID ( SLOT_2_AXI_RVALID ),
      .SLOT_2_AXI_RREADY ( SLOT_2_AXI_RREADY ),
      .SLOT_2_AXIS_ACLK ( SLOT_2_AXIS_ACLK ),
      .SLOT_2_AXIS_ARESETN ( SLOT_2_AXIS_ARESETN ),
      .SLOT_2_AXIS_TVALID ( SLOT_2_AXIS_TVALID ),
      .SLOT_2_AXIS_TREADY ( SLOT_2_AXIS_TREADY ),
      .SLOT_2_AXIS_TDATA ( SLOT_2_AXIS_TDATA ),
      .SLOT_2_AXIS_TSTRB ( SLOT_2_AXIS_TSTRB ),
      .SLOT_2_AXIS_TKEEP ( SLOT_2_AXIS_TKEEP ),
      .SLOT_2_AXIS_TLAST ( SLOT_2_AXIS_TLAST ),
      .SLOT_2_AXIS_TID ( SLOT_2_AXIS_TID ),
      .SLOT_2_AXIS_TDEST ( SLOT_2_AXIS_TDEST ),
      .SLOT_2_AXIS_TUSER ( SLOT_2_AXIS_TUSER ),
      .SLOT_3_AXI_ACLK ( SLOT_3_AXI_ACLK ),
      .SLOT_3_AXI_ARESETN ( SLOT_3_AXI_ARESETN ),
      .SLOT_3_AXI_AWID ( SLOT_3_AXI_AWID ),
      .SLOT_3_AXI_AWADDR ( SLOT_3_AXI_AWADDR ),
      .SLOT_3_AXI_AWLEN ( SLOT_3_AXI_AWLEN ),
      .SLOT_3_AXI_AWPROT ( SLOT_3_AXI_AWPROT ),
      .SLOT_3_AXI_AWSIZE ( SLOT_3_AXI_AWSIZE ),
      .SLOT_3_AXI_AWBURST ( SLOT_3_AXI_AWBURST ),
      .SLOT_3_AXI_AWCACHE ( SLOT_3_AXI_AWCACHE ),
      .SLOT_3_AXI_AWLOCK ( SLOT_3_AXI_AWLOCK ),
      .SLOT_3_AXI_AWVALID ( SLOT_3_AXI_AWVALID ),
      .SLOT_3_AXI_AWREADY ( SLOT_3_AXI_AWREADY ),
      .SLOT_3_AXI_WDATA ( SLOT_3_AXI_WDATA ),
      .SLOT_3_AXI_WSTRB ( SLOT_3_AXI_WSTRB ),
      .SLOT_3_AXI_WLAST ( SLOT_3_AXI_WLAST ),
      .SLOT_3_AXI_WVALID ( SLOT_3_AXI_WVALID ),
      .SLOT_3_AXI_WREADY ( SLOT_3_AXI_WREADY ),
      .SLOT_3_AXI_BID ( SLOT_3_AXI_BID ),
      .SLOT_3_AXI_BRESP ( SLOT_3_AXI_BRESP ),
      .SLOT_3_AXI_BVALID ( SLOT_3_AXI_BVALID ),
      .SLOT_3_AXI_BREADY ( SLOT_3_AXI_BREADY ),
      .SLOT_3_AXI_ARID ( SLOT_3_AXI_ARID ),
      .SLOT_3_AXI_ARADDR ( SLOT_3_AXI_ARADDR ),
      .SLOT_3_AXI_ARLEN ( SLOT_3_AXI_ARLEN ),
      .SLOT_3_AXI_ARSIZE ( SLOT_3_AXI_ARSIZE ),
      .SLOT_3_AXI_ARBURST ( SLOT_3_AXI_ARBURST ),
      .SLOT_3_AXI_ARPROT ( SLOT_3_AXI_ARPROT ),
      .SLOT_3_AXI_ARCACHE ( SLOT_3_AXI_ARCACHE ),
      .SLOT_3_AXI_ARLOCK ( SLOT_3_AXI_ARLOCK ),
      .SLOT_3_AXI_ARVALID ( SLOT_3_AXI_ARVALID ),
      .SLOT_3_AXI_ARREADY ( SLOT_3_AXI_ARREADY ),
      .SLOT_3_AXI_RID ( SLOT_3_AXI_RID ),
      .SLOT_3_AXI_RDATA ( SLOT_3_AXI_RDATA ),
      .SLOT_3_AXI_RRESP ( SLOT_3_AXI_RRESP ),
      .SLOT_3_AXI_RLAST ( SLOT_3_AXI_RLAST ),
      .SLOT_3_AXI_RVALID ( SLOT_3_AXI_RVALID ),
      .SLOT_3_AXI_RREADY ( SLOT_3_AXI_RREADY ),
      .SLOT_3_AXIS_ACLK ( SLOT_3_AXIS_ACLK ),
      .SLOT_3_AXIS_ARESETN ( SLOT_3_AXIS_ARESETN ),
      .SLOT_3_AXIS_TVALID ( SLOT_3_AXIS_TVALID ),
      .SLOT_3_AXIS_TREADY ( SLOT_3_AXIS_TREADY ),
      .SLOT_3_AXIS_TDATA ( SLOT_3_AXIS_TDATA ),
      .SLOT_3_AXIS_TSTRB ( SLOT_3_AXIS_TSTRB ),
      .SLOT_3_AXIS_TKEEP ( SLOT_3_AXIS_TKEEP ),
      .SLOT_3_AXIS_TLAST ( SLOT_3_AXIS_TLAST ),
      .SLOT_3_AXIS_TID ( SLOT_3_AXIS_TID ),
      .SLOT_3_AXIS_TDEST ( SLOT_3_AXIS_TDEST ),
      .SLOT_3_AXIS_TUSER ( SLOT_3_AXIS_TUSER ),
      .SLOT_4_AXI_ACLK ( SLOT_4_AXI_ACLK ),
      .SLOT_4_AXI_ARESETN ( SLOT_4_AXI_ARESETN ),
      .SLOT_4_AXI_AWID ( SLOT_4_AXI_AWID ),
      .SLOT_4_AXI_AWADDR ( SLOT_4_AXI_AWADDR ),
      .SLOT_4_AXI_AWLEN ( SLOT_4_AXI_AWLEN ),
      .SLOT_4_AXI_AWPROT ( SLOT_4_AXI_AWPROT ),
      .SLOT_4_AXI_AWSIZE ( SLOT_4_AXI_AWSIZE ),
      .SLOT_4_AXI_AWBURST ( SLOT_4_AXI_AWBURST ),
      .SLOT_4_AXI_AWCACHE ( SLOT_4_AXI_AWCACHE ),
      .SLOT_4_AXI_AWLOCK ( SLOT_4_AXI_AWLOCK ),
      .SLOT_4_AXI_AWVALID ( SLOT_4_AXI_AWVALID ),
      .SLOT_4_AXI_AWREADY ( SLOT_4_AXI_AWREADY ),
      .SLOT_4_AXI_WDATA ( SLOT_4_AXI_WDATA ),
      .SLOT_4_AXI_WSTRB ( SLOT_4_AXI_WSTRB ),
      .SLOT_4_AXI_WLAST ( SLOT_4_AXI_WLAST ),
      .SLOT_4_AXI_WVALID ( SLOT_4_AXI_WVALID ),
      .SLOT_4_AXI_WREADY ( SLOT_4_AXI_WREADY ),
      .SLOT_4_AXI_BID ( SLOT_4_AXI_BID ),
      .SLOT_4_AXI_BRESP ( SLOT_4_AXI_BRESP ),
      .SLOT_4_AXI_BVALID ( SLOT_4_AXI_BVALID ),
      .SLOT_4_AXI_BREADY ( SLOT_4_AXI_BREADY ),
      .SLOT_4_AXI_ARID ( SLOT_4_AXI_ARID ),
      .SLOT_4_AXI_ARADDR ( SLOT_4_AXI_ARADDR ),
      .SLOT_4_AXI_ARLEN ( SLOT_4_AXI_ARLEN ),
      .SLOT_4_AXI_ARSIZE ( SLOT_4_AXI_ARSIZE ),
      .SLOT_4_AXI_ARBURST ( SLOT_4_AXI_ARBURST ),
      .SLOT_4_AXI_ARPROT ( SLOT_4_AXI_ARPROT ),
      .SLOT_4_AXI_ARCACHE ( SLOT_4_AXI_ARCACHE ),
      .SLOT_4_AXI_ARLOCK ( SLOT_4_AXI_ARLOCK ),
      .SLOT_4_AXI_ARVALID ( SLOT_4_AXI_ARVALID ),
      .SLOT_4_AXI_ARREADY ( SLOT_4_AXI_ARREADY ),
      .SLOT_4_AXI_RID ( SLOT_4_AXI_RID ),
      .SLOT_4_AXI_RDATA ( SLOT_4_AXI_RDATA ),
      .SLOT_4_AXI_RRESP ( SLOT_4_AXI_RRESP ),
      .SLOT_4_AXI_RLAST ( SLOT_4_AXI_RLAST ),
      .SLOT_4_AXI_RVALID ( SLOT_4_AXI_RVALID ),
      .SLOT_4_AXI_RREADY ( SLOT_4_AXI_RREADY ),
      .SLOT_4_AXIS_ACLK ( SLOT_4_AXIS_ACLK ),
      .SLOT_4_AXIS_ARESETN ( SLOT_4_AXIS_ARESETN ),
      .SLOT_4_AXIS_TVALID ( SLOT_4_AXIS_TVALID ),
      .SLOT_4_AXIS_TREADY ( SLOT_4_AXIS_TREADY ),
      .SLOT_4_AXIS_TDATA ( SLOT_4_AXIS_TDATA ),
      .SLOT_4_AXIS_TSTRB ( SLOT_4_AXIS_TSTRB ),
      .SLOT_4_AXIS_TKEEP ( SLOT_4_AXIS_TKEEP ),
      .SLOT_4_AXIS_TLAST ( SLOT_4_AXIS_TLAST ),
      .SLOT_4_AXIS_TID ( SLOT_4_AXIS_TID ),
      .SLOT_4_AXIS_TDEST ( SLOT_4_AXIS_TDEST ),
      .SLOT_4_AXIS_TUSER ( SLOT_4_AXIS_TUSER ),
      .SLOT_5_AXI_ACLK ( SLOT_5_AXI_ACLK ),
      .SLOT_5_AXI_ARESETN ( SLOT_5_AXI_ARESETN ),
      .SLOT_5_AXI_AWID ( SLOT_5_AXI_AWID ),
      .SLOT_5_AXI_AWADDR ( SLOT_5_AXI_AWADDR ),
      .SLOT_5_AXI_AWLEN ( SLOT_5_AXI_AWLEN ),
      .SLOT_5_AXI_AWPROT ( SLOT_5_AXI_AWPROT ),
      .SLOT_5_AXI_AWSIZE ( SLOT_5_AXI_AWSIZE ),
      .SLOT_5_AXI_AWBURST ( SLOT_5_AXI_AWBURST ),
      .SLOT_5_AXI_AWCACHE ( SLOT_5_AXI_AWCACHE ),
      .SLOT_5_AXI_AWLOCK ( SLOT_5_AXI_AWLOCK ),
      .SLOT_5_AXI_AWVALID ( SLOT_5_AXI_AWVALID ),
      .SLOT_5_AXI_AWREADY ( SLOT_5_AXI_AWREADY ),
      .SLOT_5_AXI_WDATA ( SLOT_5_AXI_WDATA ),
      .SLOT_5_AXI_WSTRB ( SLOT_5_AXI_WSTRB ),
      .SLOT_5_AXI_WLAST ( SLOT_5_AXI_WLAST ),
      .SLOT_5_AXI_WVALID ( SLOT_5_AXI_WVALID ),
      .SLOT_5_AXI_WREADY ( SLOT_5_AXI_WREADY ),
      .SLOT_5_AXI_BID ( SLOT_5_AXI_BID ),
      .SLOT_5_AXI_BRESP ( SLOT_5_AXI_BRESP ),
      .SLOT_5_AXI_BVALID ( SLOT_5_AXI_BVALID ),
      .SLOT_5_AXI_BREADY ( SLOT_5_AXI_BREADY ),
      .SLOT_5_AXI_ARID ( SLOT_5_AXI_ARID ),
      .SLOT_5_AXI_ARADDR ( SLOT_5_AXI_ARADDR ),
      .SLOT_5_AXI_ARLEN ( SLOT_5_AXI_ARLEN ),
      .SLOT_5_AXI_ARSIZE ( SLOT_5_AXI_ARSIZE ),
      .SLOT_5_AXI_ARBURST ( SLOT_5_AXI_ARBURST ),
      .SLOT_5_AXI_ARPROT ( SLOT_5_AXI_ARPROT ),
      .SLOT_5_AXI_ARCACHE ( SLOT_5_AXI_ARCACHE ),
      .SLOT_5_AXI_ARLOCK ( SLOT_5_AXI_ARLOCK ),
      .SLOT_5_AXI_ARVALID ( SLOT_5_AXI_ARVALID ),
      .SLOT_5_AXI_ARREADY ( SLOT_5_AXI_ARREADY ),
      .SLOT_5_AXI_RID ( SLOT_5_AXI_RID ),
      .SLOT_5_AXI_RDATA ( SLOT_5_AXI_RDATA ),
      .SLOT_5_AXI_RRESP ( SLOT_5_AXI_RRESP ),
      .SLOT_5_AXI_RLAST ( SLOT_5_AXI_RLAST ),
      .SLOT_5_AXI_RVALID ( SLOT_5_AXI_RVALID ),
      .SLOT_5_AXI_RREADY ( SLOT_5_AXI_RREADY ),
      .SLOT_5_AXIS_ACLK ( SLOT_5_AXIS_ACLK ),
      .SLOT_5_AXIS_ARESETN ( SLOT_5_AXIS_ARESETN ),
      .SLOT_5_AXIS_TVALID ( SLOT_5_AXIS_TVALID ),
      .SLOT_5_AXIS_TREADY ( SLOT_5_AXIS_TREADY ),
      .SLOT_5_AXIS_TDATA ( SLOT_5_AXIS_TDATA ),
      .SLOT_5_AXIS_TSTRB ( SLOT_5_AXIS_TSTRB ),
      .SLOT_5_AXIS_TKEEP ( SLOT_5_AXIS_TKEEP ),
      .SLOT_5_AXIS_TLAST ( SLOT_5_AXIS_TLAST ),
      .SLOT_5_AXIS_TID ( SLOT_5_AXIS_TID ),
      .SLOT_5_AXIS_TDEST ( SLOT_5_AXIS_TDEST ),
      .SLOT_5_AXIS_TUSER ( SLOT_5_AXIS_TUSER ),
      .SLOT_6_AXI_ACLK ( SLOT_6_AXI_ACLK ),
      .SLOT_6_AXI_ARESETN ( SLOT_6_AXI_ARESETN ),
      .SLOT_6_AXI_AWID ( SLOT_6_AXI_AWID ),
      .SLOT_6_AXI_AWADDR ( SLOT_6_AXI_AWADDR ),
      .SLOT_6_AXI_AWLEN ( SLOT_6_AXI_AWLEN ),
      .SLOT_6_AXI_AWPROT ( SLOT_6_AXI_AWPROT ),
      .SLOT_6_AXI_AWSIZE ( SLOT_6_AXI_AWSIZE ),
      .SLOT_6_AXI_AWBURST ( SLOT_6_AXI_AWBURST ),
      .SLOT_6_AXI_AWCACHE ( SLOT_6_AXI_AWCACHE ),
      .SLOT_6_AXI_AWLOCK ( SLOT_6_AXI_AWLOCK ),
      .SLOT_6_AXI_AWVALID ( SLOT_6_AXI_AWVALID ),
      .SLOT_6_AXI_AWREADY ( SLOT_6_AXI_AWREADY ),
      .SLOT_6_AXI_WDATA ( SLOT_6_AXI_WDATA ),
      .SLOT_6_AXI_WSTRB ( SLOT_6_AXI_WSTRB ),
      .SLOT_6_AXI_WLAST ( SLOT_6_AXI_WLAST ),
      .SLOT_6_AXI_WVALID ( SLOT_6_AXI_WVALID ),
      .SLOT_6_AXI_WREADY ( SLOT_6_AXI_WREADY ),
      .SLOT_6_AXI_BID ( SLOT_6_AXI_BID ),
      .SLOT_6_AXI_BRESP ( SLOT_6_AXI_BRESP ),
      .SLOT_6_AXI_BVALID ( SLOT_6_AXI_BVALID ),
      .SLOT_6_AXI_BREADY ( SLOT_6_AXI_BREADY ),
      .SLOT_6_AXI_ARID ( SLOT_6_AXI_ARID ),
      .SLOT_6_AXI_ARADDR ( SLOT_6_AXI_ARADDR ),
      .SLOT_6_AXI_ARLEN ( SLOT_6_AXI_ARLEN ),
      .SLOT_6_AXI_ARSIZE ( SLOT_6_AXI_ARSIZE ),
      .SLOT_6_AXI_ARBURST ( SLOT_6_AXI_ARBURST ),
      .SLOT_6_AXI_ARPROT ( SLOT_6_AXI_ARPROT ),
      .SLOT_6_AXI_ARCACHE ( SLOT_6_AXI_ARCACHE ),
      .SLOT_6_AXI_ARLOCK ( SLOT_6_AXI_ARLOCK ),
      .SLOT_6_AXI_ARVALID ( SLOT_6_AXI_ARVALID ),
      .SLOT_6_AXI_ARREADY ( SLOT_6_AXI_ARREADY ),
      .SLOT_6_AXI_RID ( SLOT_6_AXI_RID ),
      .SLOT_6_AXI_RDATA ( SLOT_6_AXI_RDATA ),
      .SLOT_6_AXI_RRESP ( SLOT_6_AXI_RRESP ),
      .SLOT_6_AXI_RLAST ( SLOT_6_AXI_RLAST ),
      .SLOT_6_AXI_RVALID ( SLOT_6_AXI_RVALID ),
      .SLOT_6_AXI_RREADY ( SLOT_6_AXI_RREADY ),
      .SLOT_6_AXIS_ACLK ( SLOT_6_AXIS_ACLK ),
      .SLOT_6_AXIS_ARESETN ( SLOT_6_AXIS_ARESETN ),
      .SLOT_6_AXIS_TVALID ( SLOT_6_AXIS_TVALID ),
      .SLOT_6_AXIS_TREADY ( SLOT_6_AXIS_TREADY ),
      .SLOT_6_AXIS_TDATA ( SLOT_6_AXIS_TDATA ),
      .SLOT_6_AXIS_TSTRB ( SLOT_6_AXIS_TSTRB ),
      .SLOT_6_AXIS_TKEEP ( SLOT_6_AXIS_TKEEP ),
      .SLOT_6_AXIS_TLAST ( SLOT_6_AXIS_TLAST ),
      .SLOT_6_AXIS_TID ( SLOT_6_AXIS_TID ),
      .SLOT_6_AXIS_TDEST ( SLOT_6_AXIS_TDEST ),
      .SLOT_6_AXIS_TUSER ( SLOT_6_AXIS_TUSER ),
      .SLOT_7_AXI_ACLK ( SLOT_7_AXI_ACLK ),
      .SLOT_7_AXI_ARESETN ( SLOT_7_AXI_ARESETN ),
      .SLOT_7_AXI_AWID ( SLOT_7_AXI_AWID ),
      .SLOT_7_AXI_AWADDR ( SLOT_7_AXI_AWADDR ),
      .SLOT_7_AXI_AWLEN ( SLOT_7_AXI_AWLEN ),
      .SLOT_7_AXI_AWPROT ( SLOT_7_AXI_AWPROT ),
      .SLOT_7_AXI_AWSIZE ( SLOT_7_AXI_AWSIZE ),
      .SLOT_7_AXI_AWBURST ( SLOT_7_AXI_AWBURST ),
      .SLOT_7_AXI_AWCACHE ( SLOT_7_AXI_AWCACHE ),
      .SLOT_7_AXI_AWLOCK ( SLOT_7_AXI_AWLOCK ),
      .SLOT_7_AXI_AWVALID ( SLOT_7_AXI_AWVALID ),
      .SLOT_7_AXI_AWREADY ( SLOT_7_AXI_AWREADY ),
      .SLOT_7_AXI_WDATA ( SLOT_7_AXI_WDATA ),
      .SLOT_7_AXI_WSTRB ( SLOT_7_AXI_WSTRB ),
      .SLOT_7_AXI_WLAST ( SLOT_7_AXI_WLAST ),
      .SLOT_7_AXI_WVALID ( SLOT_7_AXI_WVALID ),
      .SLOT_7_AXI_WREADY ( SLOT_7_AXI_WREADY ),
      .SLOT_7_AXI_BID ( SLOT_7_AXI_BID ),
      .SLOT_7_AXI_BRESP ( SLOT_7_AXI_BRESP ),
      .SLOT_7_AXI_BVALID ( SLOT_7_AXI_BVALID ),
      .SLOT_7_AXI_BREADY ( SLOT_7_AXI_BREADY ),
      .SLOT_7_AXI_ARID ( SLOT_7_AXI_ARID ),
      .SLOT_7_AXI_ARADDR ( SLOT_7_AXI_ARADDR ),
      .SLOT_7_AXI_ARLEN ( SLOT_7_AXI_ARLEN ),
      .SLOT_7_AXI_ARSIZE ( SLOT_7_AXI_ARSIZE ),
      .SLOT_7_AXI_ARBURST ( SLOT_7_AXI_ARBURST ),
      .SLOT_7_AXI_ARPROT ( SLOT_7_AXI_ARPROT ),
      .SLOT_7_AXI_ARCACHE ( SLOT_7_AXI_ARCACHE ),
      .SLOT_7_AXI_ARLOCK ( SLOT_7_AXI_ARLOCK ),
      .SLOT_7_AXI_ARVALID ( SLOT_7_AXI_ARVALID ),
      .SLOT_7_AXI_ARREADY ( SLOT_7_AXI_ARREADY ),
      .SLOT_7_AXI_RID ( SLOT_7_AXI_RID ),
      .SLOT_7_AXI_RDATA ( SLOT_7_AXI_RDATA ),
      .SLOT_7_AXI_RRESP ( SLOT_7_AXI_RRESP ),
      .SLOT_7_AXI_RLAST ( SLOT_7_AXI_RLAST ),
      .SLOT_7_AXI_RVALID ( SLOT_7_AXI_RVALID ),
      .SLOT_7_AXI_RREADY ( SLOT_7_AXI_RREADY ),
      .SLOT_7_AXIS_ACLK ( SLOT_7_AXIS_ACLK ),
      .SLOT_7_AXIS_ARESETN ( SLOT_7_AXIS_ARESETN ),
      .SLOT_7_AXIS_TVALID ( SLOT_7_AXIS_TVALID ),
      .SLOT_7_AXIS_TREADY ( SLOT_7_AXIS_TREADY ),
      .SLOT_7_AXIS_TDATA ( SLOT_7_AXIS_TDATA ),
      .SLOT_7_AXIS_TSTRB ( SLOT_7_AXIS_TSTRB ),
      .SLOT_7_AXIS_TKEEP ( SLOT_7_AXIS_TKEEP ),
      .SLOT_7_AXIS_TLAST ( SLOT_7_AXIS_TLAST ),
      .SLOT_7_AXIS_TID ( SLOT_7_AXIS_TID ),
      .SLOT_7_AXIS_TDEST ( SLOT_7_AXIS_TDEST ),
      .SLOT_7_AXIS_TUSER ( SLOT_7_AXIS_TUSER ),
      .EXT_CLK_0 ( EXT_CLK_0 ),
      .EXT_RSTN_0 ( EXT_RSTN_0 ),
      .EXT_EVENT_0_CNT_START ( EXT_EVENT_0_CNT_START ),
      .EXT_EVENT_0_CNT_STOP ( EXT_EVENT_0_CNT_STOP ),
      .EXT_EVENT_0 ( EXT_EVENT_0 ),
      .EXT_CLK_1 ( EXT_CLK_1 ),
      .EXT_RSTN_1 ( EXT_RSTN_1 ),
      .EXT_EVENT_1_CNT_START ( EXT_EVENT_1_CNT_START ),
      .EXT_EVENT_1_CNT_STOP ( EXT_EVENT_1_CNT_STOP ),
      .EXT_EVENT_1 ( EXT_EVENT_1 ),
      .EXT_CLK_2 ( EXT_CLK_2 ),
      .EXT_RSTN_2 ( EXT_RSTN_2 ),
      .EXT_EVENT_2_CNT_START ( EXT_EVENT_2_CNT_START ),
      .EXT_EVENT_2_CNT_STOP ( EXT_EVENT_2_CNT_STOP ),
      .EXT_EVENT_2 ( EXT_EVENT_2 ),
      .EXT_CLK_3 ( EXT_CLK_3 ),
      .EXT_RSTN_3 ( EXT_RSTN_3 ),
      .EXT_EVENT_3_CNT_START ( EXT_EVENT_3_CNT_START ),
      .EXT_EVENT_3_CNT_STOP ( EXT_EVENT_3_CNT_STOP ),
      .EXT_EVENT_3 ( EXT_EVENT_3 ),
      .EXT_CLK_4 ( EXT_CLK_4 ),
      .EXT_RSTN_4 ( EXT_RSTN_4 ),
      .EXT_EVENT_4_CNT_START ( EXT_EVENT_4_CNT_START ),
      .EXT_EVENT_4_CNT_STOP ( EXT_EVENT_4_CNT_STOP ),
      .EXT_EVENT_4 ( EXT_EVENT_4 ),
      .EXT_CLK_5 ( EXT_CLK_5 ),
      .EXT_RSTN_5 ( EXT_RSTN_5 ),
      .EXT_EVENT_5_CNT_START ( EXT_EVENT_5_CNT_START ),
      .EXT_EVENT_5_CNT_STOP ( EXT_EVENT_5_CNT_STOP ),
      .EXT_EVENT_5 ( EXT_EVENT_5 ),
      .EXT_CLK_6 ( EXT_CLK_6 ),
      .EXT_RSTN_6 ( EXT_RSTN_6 ),
      .EXT_EVENT_6_CNT_START ( EXT_EVENT_6_CNT_START ),
      .EXT_EVENT_6_CNT_STOP ( EXT_EVENT_6_CNT_STOP ),
      .EXT_EVENT_6 ( EXT_EVENT_6 ),
      .EXT_CLK_7 ( EXT_CLK_7 ),
      .EXT_RSTN_7 ( EXT_RSTN_7 ),
      .EXT_EVENT_7_CNT_START ( EXT_EVENT_7_CNT_START ),
      .EXT_EVENT_7_CNT_STOP ( EXT_EVENT_7_CNT_STOP ),
      .EXT_EVENT_7 ( EXT_EVENT_7 ),
      .SLOT_0_EXT_TRIG ( SLOT_0_EXT_TRIG ),
      .SLOT_1_EXT_TRIG ( SLOT_1_EXT_TRIG ),
      .SLOT_2_EXT_TRIG ( SLOT_2_EXT_TRIG ),
      .SLOT_3_EXT_TRIG ( SLOT_3_EXT_TRIG ),
      .SLOT_4_EXT_TRIG ( SLOT_4_EXT_TRIG ),
      .SLOT_5_EXT_TRIG ( SLOT_5_EXT_TRIG ),
      .SLOT_6_EXT_TRIG ( SLOT_6_EXT_TRIG ),
      .SLOT_7_EXT_TRIG ( SLOT_7_EXT_TRIG ),
      .CAPTURE_EVENT ( CAPTURE_EVENT ),
      .RESET_EVENT ( RESET_EVENT ),
      .M_AXIS_ACLK ( M_AXIS_ACLK ),
      .M_AXIS_ARESETN ( M_AXIS_ARESETN ),
      .M_AXIS_TDATA ( M_AXIS_TDATA ),
      .M_AXIS_TSTRB ( M_AXIS_TSTRB ),
      .M_AXIS_TVALID ( M_AXIS_TVALID ),
      .M_AXIS_TID ( M_AXIS_TID ),
      .M_AXIS_TREADY ( M_AXIS_TREADY ),
      .CORE_ACLK ( CORE_ACLK ),
      .CORE_ARESETN ( CORE_ARESETN ),
      .INTERRUPT ( INTERRUPT )
    );

endmodule

